module enemy_mgr (
    input  wire clk,
    input  wire rst
);

endmodule //enemy_mgr